library verilog;
use verilog.vl_types.all;
entity out_FSM_vlg_vec_tst is
end out_FSM_vlg_vec_tst;
