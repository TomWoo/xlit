module output_FSM(
input clk,
input rst,
input [63:0] frame_count
//input []
);



endmodule
