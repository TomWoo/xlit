library verilog;
use verilog.vl_types.all;
entity xmitTop_vlg_vec_tst is
end xmitTop_vlg_vec_tst;
