library ieee;
use ieee.std_logic_1164.all;

entity in_FSM is 
port(
	in_frame:				in std_logic_vector(7 downto 0);
	in_priority:			in std_logic;
	in_low_overflow:		in std_logic;
	in_hi_overflow:		in std_logic;
	in_f_rdv:				in std_logic;
	out_m_discard_en:		out std_logic;
	--out_m_discard_frame:	out std_logic_vector(7 downto 0);
	out_frame:				out std_logic_vector(7 downto 0);
	out_wren:				out std_logic;
	out_priority: 			out std_logic;
	clk_sys:					in std_logic;
	reset:					in std_logic			
);
end in_FSM;

architecture arch of in_FSM is
	type numstate is (start_state, frame_state, end_state);
	
begin

	process(clk_sys, reset)
	begin
		if(reset = '1') then
			out_m_discard_en <= '0';
		elsif (clk_sys'event and clk_sys='1') then
			if ((in_low_overflow = '1' and in_priority='0') or (in_hi_overflow='1' and in_priority='1')) then
				out_m_discard_en <= '1';
			else
				out_m_discard_en <= '0';
			end if;
		end if;
	end process;
	
	process(clk_sys, reset)
	begin
		if(reset = '1') then
			out_wren <= '0';
		elsif (clk_sys'event and clk_sys='1') then
			out_wren <= in_f_rdv;
		end if;
	end process;
	
	process(clk_sys, reset) begin
		out_frame <= in_frame;
		out_priority <= in_priority;
	end process;
	/*
	process(clk_sys, reset) begin
		if(reset = '1') then
			
		end if;
	end process;
	*/
end arch;
