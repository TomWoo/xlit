library verilog;
use verilog.vl_types.all;
entity in_FSM_vlg_vec_tst is
end in_FSM_vlg_vec_tst;
